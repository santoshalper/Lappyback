example lowpass
.model DMOD D(vj=1.7)
r1 1 2 2.2k
df 2 0 DMOD
dr 0 2 DMOD
c2 2 0 .1u
v1 1 0 pulse(0 5 0 1.14m 1.14m 0 2.28m)
r2 2 0 100k
*v2 1 0 dc 0 ac 2.5
.option noacct
*.ac oct 10 20 20k
.tran 1ms 10ms
.end
